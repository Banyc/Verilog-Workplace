`ifndef __Alu32b_simple_enumAluOp_vh__
`define __Alu32b_simple_enumAluOp_vh__

`define Alu32b_simple_aluOp_and 4'b0000
`define Alu32b_simple_aluOp_or  4'b0001
`define Alu32b_simple_aluOp_add 4'b0010
`define Alu32b_simple_aluOp_sub 4'b0110
`define Alu32b_simple_aluOp_slt 4'b0111
`define Alu32b_simple_aluOp_nor 4'b1100

`endif
