
`include "./Components/multiplier/Divider32b.v"

module Top(
    
);

endmodule // Top
