`ifndef __EnumFunct7_vh__
`define __EnumFunct7_vh__

// riscv-spec.pdf #130

`define riscv32_funct7_SLLI  7'b0000000
`define riscv32_funct7_SRLI  7'b0000000
`define riscv32_funct7_SRAI  7'b0100000
`define riscv32_funct7_ADD   7'b0000000
`define riscv32_funct7_SUB   7'b0100000
`define riscv32_funct7_SLL   7'b0000000
`define riscv32_funct7_SLT   7'b0000000
`define riscv32_funct7_SLTU  7'b0000000
`define riscv32_funct7_XOR   7'b0000000
`define riscv32_funct7_SRL   7'b0000000
`define riscv32_funct7_SRA   7'b0100000
`define riscv32_funct7_OR    7'b0000000
`define riscv32_funct7_AND   7'b0000000

`endif
