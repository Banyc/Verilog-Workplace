`ifndef __Alu32b_extended_enumAluOp_vh__
`define __Alu32b_extended_enumAluOp_vh__

`define Alu32b_extended_aluOp_and  4'b0000
`define Alu32b_extended_aluOp_or   4'b0001
`define Alu32b_extended_aluOp_add  4'b0010
`define Alu32b_extended_aluOp_sub  4'b0110
`define Alu32b_extended_aluOp_slt  4'b0111
`define Alu32b_extended_aluOp_nor  4'b1100

`define Alu32b_extended_aluOp_sll  4'b1011
`define Alu32b_extended_aluOp_srl  4'b1111
`define Alu32b_extended_aluOp_sra  4'b1010
`define Alu32b_extended_aluOp_xor  4'b1110
`define Alu32b_extended_aluOp_sltu 4'b1000

`endif
