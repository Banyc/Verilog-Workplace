`ifndef __EnumInstructionTypes_vh__
`define __EnumInstructionTypes_vh__

`define riscv_instructionType_R   0
`define riscv_instructionType_I   1
`define riscv_instructionType_S   2
`define riscv_instructionType_SB  3
`define riscv_instructionType_U   4
`define riscv_instructionType_UJ  5
`define riscv_instructionType_undefined  6

`endif
